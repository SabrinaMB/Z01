library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Nor8Way is
	port ( 
			a:   in  STD_LOGIC;
			b:   in  STD_LOGIC;
			c:   in  STD_LOGIC;
			d:   in  STD_LOGIC;
			e:   in  STD_LOGIC;
			f:   in  STD_LOGIC;
			g:   in  STD_LOGIC;
			h:   in  STD_LOGIC;
			q:   out STD_LOGIC);
<<<<<<< HEAD
end Nor8Way;

architecture n8 of Nor8Way is
begin
	q <= not (a or b or c or d or e or f or g or h);
end n8;
=======
end entity;
>>>>>>> upstream/master
