-- Elementos de Sistemas
-- by Phelipe Muller
-- Register32.vhd

Library ieee;
use ieee.std_logic_1164.all;

-- by Luciano Soares
-- Register32.vhd

Library ieee; 
use ieee.std_logic_1164.all;
  
entity Register32 is
	port(
		clock:   in STD_LOGIC;
		input:   in STD_LOGIC_VECTOR(31 downto 0);
		load:    in STD_LOGIC;
		output: out STD_LOGIC_VECTOR(31 downto 0)
	);
end entity;


architecture arch of Register32 is

  component Register16 is
    port(
    clock:   in STD_LOGIC;
		input:   in STD_LOGIC_VECTOR(15 downto 0);
		load:    in STD_LOGIC;
		output: out STD_LOGIC_VECTOR(15 downto 0)
	);
  end component;

begin
  R1 : Register16 PORT MAP(clock,input(15 downto 0),load,output(15 downto 0));
  R2 : Register16 PORT MAP(clock,input(31 downto 16),load,output(31 downto 16));

end architecture;

