library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity DMux2Way is
	port ( 
			a:   in  STD_LOGIC;
			sel: in  STD_LOGIC;
			q0:  out STD_LOGIC;
			q1:  out STD_LOGIC);
<<<<<<< HEAD
end entity;

architecture this_DMux of DMux2Way is
begin

   q1 <= a when(sel = '1') else '0';
   q0 <= a when(sel = '0') else '0';

end this_DMux;
=======
end entity
>>>>>>> upstream/master
