library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Not16 is
	port ( 
			a:   in  STD_LOGIC_VECTOR(15 downto 0);
			q:   out STD_LOGIC_VECTOR(15 downto 0));
<<<<<<< HEAD
end entity;

architecture this_not16 of Not16 is
begin
	q <= not a;
end this_not16;
=======
end entity;
>>>>>>> upstream/master
